
module fwspi_initiator_hdl_top;
endmodule

