`include "uvm_macros.svh"

module fwspi_initiator_hvl_top;
    import uvm_pkg::*;

    fwspi_initiator_hdl_top u_top();

endmodule
